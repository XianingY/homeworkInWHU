`define alu_add 4'b0010
`define alu_sub 4'b0110
`define alu_and 4'b0000
`define alu_or 4'b0001
`define alu_xor 4'b0011
`define alu_leftlogical 4'b0100
`define alu_rightlogical 4'b0101
`define alu_right 4'b0111
`define alu_slt 4'b1000
`define alu_sltu 4'b1001

`define alu_bne 4'b1010
`define alu_blt 4'b1011
`define alu_bge 4'b1100
`define alu_bltu 4'b1101
`define alu_bgeu 4'b1111

`define jump_bne 3'b000
`define jump_blt 3'b001
`define jump_bge 3'b010
`define jump_bltu 3'b011
`define jump_bgeu 3'b100
`define jump_beq 3'b101
`define jump_jalr 3'b110
`define jump_jal 3'b111
