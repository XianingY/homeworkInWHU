module PCadd1(
    input [31:0]PCIn,
    output [31:0]PCOut
    );
  
  assign PCOut=PCIn+1;
endmodule